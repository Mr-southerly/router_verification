module tb; 
  typedef mailbox #(string) s_mb;
  s_mb mb = new(8);

  initial begin  
	string intQ[$];
  end
endmodule
